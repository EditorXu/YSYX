module myseg(
	input [3:0] x,
	input en,
	output reg [7:0] HEX0
);

	reg [15:0] y;

	always@(*)
	begin
		case(y)
		16'b0000000000000001 : HEX0 = 8'b00000010;
		16'b0000000000000010 : HEX0 = 8'b10011110;
		16'b0000000000000100 : HEX0 = 8'b00100100;
		16'b0000000000001000 : HEX0 = 8'b00001100;
		16'b0000000000010000 : HEX0 = 8'b10011000;
		16'b0000000000100000 : HEX0 = 8'b01001000;
		16'b0000000001000000 : HEX0 = 8'b01000000;
		16'b0000000010000000 : HEX0 = 8'b00011110;
		16'b0000000100000000 : HEX0 = 8'b00000000;
		16'b0000001000000000 : HEX0 = 8'b00001000;
		16'b0000010000000000 : HEX0 = 8'b00010000;
		16'b0000100000000000 : HEX0 = 8'b11000000;
		16'b0001000000000000 : HEX0 = 8'b01100010;
		16'b0010000000000000 : HEX0 = 8'b10000100;
		16'b0100000000000000 : HEX0 = 8'b01100000;
		16'b1000000000000000 : HEX0 = 8'b01110000;
		default							 : HEX0 = 8'b11111111;
		endcase
	end

decode4_16 i_decode4_16(
	.x		(x),
	.en		(en),
	.y		(y)
);

endmodule 

